`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////
// Institution:     RWTH Aachen - DSP chair
// Author:          Martin Lastovka : martin.lastovka@dsp.rwth-aachen.de
// Module Name:     regmap_pckg
// Project Name:    Efficient FPGA CNN implementation
// Description:     package defining the params of the regmap (not the autogenerated register fields)
// Synthesizable:   No
///////////////////////////////////////////////////////////////////////////////////////////////


interface regmap_rd_if //interface for internal reading of the register map
#(
    parameter ADDR_WDT,
    parameter DATA_WDT
);
logic [ADDR_WDT-1:0]  rd_addr;
logic                 rd_en;
logic [DATA_WDT-1:0]  rd_data;
logic                 rd_val;

modport regmap
(
    input  rd_addr,
    input  rd_en,
    output rd_data,
    output rd_val
);

modport requester
(
    output rd_addr,
    output rd_en,
    input  rd_data,
    input  rd_val
);
endinterface

interface regmap_wr_if //interface for internal writing to the register map
#(
    parameter ADDR_WDT,
    parameter DATA_WDT
);
logic [ADDR_WDT-1:0]   wr_addr;
logic                  wr_en;
logic [DATA_WDT-1:0]   wr_data;
logic [DATA_WDT/8-1:0] wr_strb;

modport regmap
(
    input  wr_addr,
    input  wr_en,
    input  wr_data,
    input  wr_strb
);

modport requester
(
    output wr_addr,
    output wr_en,
    output wr_data,
    output wr_strb
);
endinterface

package regmap_pckg;
import regmap_reg_pckg::*;

//autogenerate with python script

//register implemented region
parameter C_REGMAP_REG_START_ADDR = C_CTRL_REG_ADDR;
parameter C_REGMAP_REG_END_ADDR = C_PERF_CACHE_STALL_UH_REG_ADDR;
parameter C_REGMAP_REG_ADDR_WDT = $clog2(C_REGMAP_REG_END_ADDR - C_REGMAP_REG_START_ADDR + 1); 
parameter C_REGMAP_REG_INT_ADDR_WDT = C_REGMAP_REG_ADDR_WDT - 2; 
parameter C_REGMAP_REG_INT_SIZE = 2**C_REGMAP_REG_INT_ADDR_WDT; 

//RAM implemented region - tensor trans. spec.
parameter C_REGMAP_TENS_TRANS_SEQ_MAX_LEN = 2**10;
parameter C_TENS_TRANS_SEQ_CNT_WDT = $clog2(C_REGMAP_TENS_TRANS_SEQ_MAX_LEN);
parameter C_REGMAP_TENS_TRANS_SPEC_WORD_CNT = (C_TENS_TRANS_CONV_DIMS_RES_1_REG_ADDR - C_TENS_TRANS_CFG_REG_ADDR)/4 + 1;

parameter C_REGMAP_RAM_START_ADDR = C_TENS_TRANS_CFG_REG_ADDR;
parameter C_REGMAP_RAM_END_ADDR = C_REGMAP_RAM_START_ADDR + 4*C_REGMAP_TENS_TRANS_SEQ_MAX_LEN*C_REGMAP_TENS_TRANS_SPEC_WORD_CNT;
parameter C_REGMAP_RAM_ADDR_WDT = $clog2(C_REGMAP_RAM_END_ADDR - C_REGMAP_RAM_START_ADDR + 1);
parameter C_REGMAP_RAM_INT_ADDR_WDT = C_REGMAP_RAM_ADDR_WDT - 2; 
parameter C_REGMAP_RAM_INT_SIZE = 2**C_REGMAP_RAM_INT_ADDR_WDT; 

parameter C_REGMAP_ADDR_WDT = $clog2(C_REGMAP_RAM_END_ADDR - C_REGMAP_REG_START_ADDR + 1); 
parameter C_REGMAP_INT_ADDR_WDT = C_REGMAP_ADDR_WDT - 2; 
parameter C_REGMAP_DATA_WDT = CSR_DATA_WIDTH;
parameter C_REGMAP_STRB_WDT = C_REGMAP_DATA_WDT/8;

endpackage